module testbench(output logic[7:0] opcode1, opcode2);